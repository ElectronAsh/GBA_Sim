`default_nettype none
`include "../gba_core_defines.vh"
`include "../gba_mmio_defines.vh"


module dma_fsm
  (input  logic mem_wait, dma_repeat,  
   input  logic enable, start,
   input  logic new_transfer, preempted,
   input  logic genIRQ,
   input  logic allowed_to_begin, xferDone,
   output logic loadCNT, loadSAD, loadDAD, stepSRC, stepDEST, storeRData,
   output logic active, write, disable_dma, set_wdata,
   output logic irq, others_cant_preempt,
   output logic reload_xfers,
   input  logic clk, rst_b);

  enum logic [2:0] {OFF, IDLE, QUEUED, READ, WRITE, PREEMPTEDREAD} cs, ns;

  always_ff @(posedge clk, negedge rst_b) begin
    if(~rst_b)
      cs <= OFF;
    else
      cs <= ns;
  end

  always_comb begin
    set_wdata = 1'b0;
    loadCNT = 1'b0;
    loadSAD = 1'b0;
    loadDAD = 1'b0;
    stepSRC = 1'b0;
    stepDEST = 1'b0;
    storeRData = 1'b0;
    active = 1'b0;
    write = 1'b0;
    disable_dma = 1'b0;
    irq = 1'b0;
    others_cant_preempt = 1'b0;
    ns = OFF;
    reload_xfers = 0;
  
    case(cs)
      OFF: begin
        if(enable && new_transfer) begin
          loadSAD = 1'b1;
          loadDAD = 1'b1;
          loadCNT = 1'b1;
          ns = IDLE;
        end
      end
      IDLE: begin
        if(enable) begin
          if(start) begin
            if(preempted || mem_wait) begin //start & (preempted || mem_wait)
              ns = QUEUED;
            end
            else if (allowed_to_begin) begin
              ns = READ;
              active = 1'b1;
            end
            else begin
                ns = IDLE;
            end
          end
          else begin //~start
            ns = IDLE;
          end
        end
      end
      QUEUED: begin
        if(enable) begin
          if(preempted || mem_wait) begin
            ns = QUEUED;
          end
          else if (allowed_to_begin) begin
            ns = READ;
            active = 1'b1;
          end
          else begin
              ns = QUEUED;
          end
        end
      end
      READ: begin
        if(mem_wait) begin
          ns = READ;
          active = 1'b1;
        end
        else if(enable) begin
          ns = WRITE;
          others_cant_preempt = 1'b1;
          storeRData = 1'b1;
          active = 1'b1;
          stepSRC = 1'b1;
          write = 1'b1;
        end
      end
      WRITE: begin
        set_wdata = 1'b1;
        if(mem_wait) begin
          ns = WRITE;
          active = 1'b1;
        end
        else if(enable) begin
          if(xferDone & dma_repeat) begin
            ns = IDLE;
            reload_xfers = 1'b1;
            irq = genIRQ;
          end
          else if(xferDone) begin
            active = 1'b1;
            ns = OFF;
            reload_xfers = 1'b1;
            disable_dma = 1'b1;
            irq = genIRQ;
          end
          else if(preempted) begin
            active = 1'b1;
            ns = PREEMPTEDREAD;
            stepDEST = 1'b1;
          end
          else begin
            ns = READ;
            active = 1'b1;
            stepDEST = 1'b1;
          end
        end
      end
      PREEMPTEDREAD: begin
        if(enable) begin
          if(preempted || mem_wait) begin
            ns = PREEMPTEDREAD;
          end
          else if (allowed_to_begin) begin
            ns = READ;
            active = 1'b1;
          end
          else begin
              ns= PREEMPTEDREAD;
          end
        end
      end

  endcase
  end

endmodule: dma_fsm

module dma_dp
  (input  logic loadCNT, loadSAD, loadDAD,
   input  logic stepSRC, stepDEST, storeRData,
   input  logic active, write, set_wdata,
   input  logic srcGamePak, destGamePak,

   output logic xferDone, new_transfer,

   input  logic [15:0] srcAddrL, srcAddrH,
   input  logic [15:0] destAddrL, destAddrH,
   input  logic [15:0] controlL, controlH,
   input  logic sound, //Can this dma unit handle sound xfers?
   input  logic reload_xfers,

   input  logic [31:0] rdata,
   output wire  [31:0] addr, wdata,
   output wire  [1:0]  size,
   output wire         wen,

   input  logic clk, rst_b
   );

  logic [31:0] old_SAD_reg;
  logic [31:0] old_DAD_reg;
  logic [31:0] old_CTL_reg;

  logic [31:0] sAddr, dAddr;
  logic [31:0] steppedSAddr, steppedDAddr;
  logic [31:0]  nextSAddr, nextDAddr;
  logic [31:0] desiredAddr;
  logic [31:0] sAddrRaw, dAddrRaw;
  logic [31:0] data;
  logic [13:0] xfers;
  logic [13:0] wordCount;

  logic xferWord;
  logic [31:0] addrStep;
  logic [31:0] targetAddr;
  logic [1:0] sCnt, dCnt;

  logic reloadDad;
  logic sadEnable;
  logic dadEnable;
  logic [1:0] size_mem_transfer;

  assign xferWord = controlH[10];
  assign size_mem_transfer = (xferWord) ? 2'b10 : 2'b01;

  assign sAddr = {4'b0, srcGamePak & sAddrRaw[27], sAddrRaw[26:0]};
  assign dAddr = {4'b0, destGamePak & dAddrRaw[27], dAddrRaw[26:0]};

  assign sadEnable = loadSAD | stepSRC;
  assign dadEnable = loadDAD | stepDEST | (loadCNT & reloadDad);

  always_comb begin //next state logic for addresses
    reloadDad = (dCnt == 2'b11);
    addrStep = xferWord ? 32'd4 : 32'd2;
    case(sCnt)
      2'b00: steppedSAddr = sAddr + addrStep;
      2'b01: steppedSAddr = sAddr - addrStep;
      2'b10: steppedSAddr = sAddr;
      2'b11: steppedSAddr = sAddr + addrStep;
    endcase
    case(dCnt)
      2'b00: steppedDAddr = dAddr + addrStep;
      2'b01: steppedDAddr = dAddr - addrStep;
      2'b10: steppedDAddr = dAddr;
      2'b11: steppedDAddr = dAddr + addrStep;
    endcase
  end

  //Handle special dma modes
  always_comb begin
    sCnt = controlH[8:7];
    dCnt = controlH[6:5];
    targetAddr = {destAddrH, destAddrL};
    if(&controlH[13:12]) begin
      if(sound) begin
        dCnt = 2'b10;
      end
      else begin
        targetAddr = 32'h0600_0000;
      end
    end
  end

  //if writing 16 bits to upper word of an address the data
  // must be in the top word of the wdata_size
  logic [31:0] wdata_size;

  assign addr = active ? desiredAddr : {32{1'bz}};
  assign wen = active ? write : 1'bz;
  assign wdata = (active & set_wdata) ? wdata_size : {32{1'bz}};
  assign size = active ? (size_mem_transfer): {32{1'bz}};

  always_comb begin
      wdata_size = data;
      if (size_mem_transfer == 2'b01 && desiredAddr[1]==1'b1)
          wdata_size[31:16] = data[15:0];
  end

  mux_2_to_1 #(32) srcAddrMux (.i0(steppedSAddr), .i1({srcAddrH, srcAddrL}), .s(loadSAD), .y(nextSAddr));
  mux_2_to_1 #(32) destAddrMux (.i0(steppedDAddr), .i1(targetAddr), .s(loadDAD | (loadCNT & reloadDad)), .y(nextDAddr));
  mux_2_to_1 #(32) addrMux (.i0(sAddr), .i1(dAddr), .s(write), .y(desiredAddr));

  register #(32) sad(.d(nextSAddr), .q(sAddrRaw), .clk, .clear(1'b0), .enable(sadEnable), .rst_b);
  register #(32) dad(.d(nextDAddr), .q(dAddrRaw), .clk, .clear(1'b0), .enable(dadEnable), .rst_b);
  register #(32) data_reg(.d(rdata), .q(data), .clk, .clear(1'b0), .enable(storeRData), .rst_b);
  counter #(14) xferCnt (.d(14'b0), .q(xfers), .clk, .enable(stepSRC), .clear(reload_xfers), .load(1'b0), .up(1'b1), .rst_b);
  logic [13:0] words_to_transfer;
  assign words_to_transfer = (sound) ? 14'd4 : controlL[13:0];
  assign xferDone = (xfers == words_to_transfer);

  //save old SAD DAD and CNT registers
  register #(32) oldsad(.d({srcAddrH, srcAddrL}), .q(old_SAD_reg), .clk, .clear(1'b0), .enable(1'b1), .rst_b);
  register #(32) olddad(.d({destAddrH, destAddrL}), .q(old_DAD_reg), .clk, .clear(1'b0), .enable(1'b1), .rst_b);
  register #(32) oldctl(.d({controlH, controlL}), .q(old_CTL_reg), .clk, .clear(1'b0), .enable(1'b1), .rst_b);

  assign new_transfer = ((old_SAD_reg != {srcAddrH, srcAddrL}) || (old_DAD_reg != {destAddrH, destAddrL}) ||
                        (old_CTL_reg != {controlH, controlL})) ? 1'b1 : 1'b0;
endmodule: dma_dp

module dma_start
  (input  logic [15:0] controlH,
   input  logic [15:0] vcount, hcount,
   input  logic sound, sound_req, //can this dma sync with sound, and are they requesting dma
   input  logic cpu_preemptable,
   output logic start, dma_stop,
   input  logic clk, rst_b);

  logic display_sync_startable;
  logic passed_go;
  logic hold_sound;

  always_ff @(posedge clk, negedge rst_b)
    if(~rst_b)
      display_sync_startable <= 1'b0;
    else
      display_sync_startable <= passed_go;

  logic sound_req_delay;
  always_ff @(posedge clk, negedge rst_b) begin
      if(~rst_b) begin
        sound_req_delay <= 1'b0;
      end
      else if (hold_sound) begin
        sound_req_delay <= sound_req_delay; //delay by one clock cycle to shorten critical path
      end
      else begin
        sound_req_delay <= sound_req;
      end
  end

  always_comb begin
    dma_stop = 1'b0; //extra control to turn off dma repeat
    passed_go = display_sync_startable;
    hold_sound = 1'b0;
    case(controlH[13:12])
      2'b00: begin
        start = cpu_preemptable;
      end
      2'b10: begin
        start = (hcount[7:0] == 8'd240 && cpu_preemptable);
      end
      2'b01: begin
        start = (vcount[7:0] == 8'd160 && cpu_preemptable);
      end
      2'b11: begin
        if(sound) begin
          if (sound_req_delay) begin
            if(cpu_preemptable) begin
              start = 1'b1;
            end
            else begin
              start = 1'b0;
              hold_sound = 1'b1;
            end
          end
          else begin
            start = 1'b0;
            hold_sound = 1'b0;
          end
        end
        else begin
          if(vcount[7:0] == 8'd02 && display_sync_startable && cpu_preemptable) begin
            start = 1'b1;
          end
          else if(vcount[7:0] == 8'd162 && cpu_preemptable) begin
            start = 1'b0;
            dma_stop = 1'b1;
            passed_go = controlH[15]; //can start now if dma is enabled
          end
          else begin
            start = 1'b0;
          end
        end
      end
    endcase
  end

endmodule: dma_start

module dma_unit
  (input  logic [15:0] controlL, controlH,
   input  logic [15:0] srcAddrL, srcAddrH,
   input  logic [15:0] destAddrL, destAddrH,

   input  logic mem_wait, preempted,
   input  logic srcGamePak, destGamePak,
   input  logic allowed_to_begin,
   input  logic cpu_preemptable,
   output logic disable_dma,
   output logic active,
   output logic irq,
   output logic others_cant_preempt,

   input  logic [31:0] rdata,
   output wire  [31:0] addr, wdata,
   output wire  [1:0]  size,
   output wire  wen,

   input  logic [15:0] vcount, hcount,
   input  logic sound, sound_req,

   input  logic clk, rst_b
   );

  logic fsm_disable;
  logic xferDone;
  logic loadCNT, loadSAD, loadDAD;
  logic stepSRC, stepDEST;
  logic storeRData;
  logic write;

  logic dma_stop;
  logic start;
  logic set_wdata;

  logic new_transfer;
  logic reload_xfers;

  assign disable_dma = fsm_disable | dma_stop;

  dma_start starter(.controlH, .vcount, .hcount, .sound, .sound_req, .start, .dma_stop, .clk, .rst_b, .cpu_preemptable);

  dma_fsm fsm(.start, .mem_wait, .dma_repeat(controlH[9]), .preempted, .enable(controlH[15]), .xferDone,
              .genIRQ(controlH[14]), .loadCNT, .loadSAD, .loadDAD, .stepSRC, .stepDEST, .storeRData, .active,
              .write, .disable_dma(fsm_disable), .irq, .clk, .rst_b, .set_wdata, .allowed_to_begin,
              .others_cant_preempt, .new_transfer, .reload_xfers);

  dma_dp datapath(.loadCNT, .loadSAD, .loadDAD, .stepSRC, .stepDEST, .storeRData, .active, .write, .srcGamePak,
                  .destGamePak, .xferDone, .srcAddrL, .srcAddrH, .destAddrL, .destAddrH, .controlL, .controlH,
                  .sound, .rdata, .addr, .wdata, .size, .wen, .clk, .rst_b, .set_wdata, .new_transfer, .reload_xfers);

endmodule: dma_unit

module dma_top
  (
  //input  logic [31:0] registers [`NUM_IO_REGS-1:0],
  	input logic [31:0] DMA0SAD_L_REG,
	input logic [31:0] DMA0SAD_H_REG,
	input logic [31:0] DMA0DAD_L_REG,
	input logic [31:0] DMA0DAD_H_REG,
	input logic [31:0] DMA0CNT_L_REG,
	input logic [31:0] DMA0CNT_H_REG,
	input logic [31:0] DMA1SAD_L_REG,
	input logic [31:0] DMA1SAD_H_REG,
	input logic [31:0] DMA1DAD_L_REG,
	input logic [31:0] DMA1DAD_H_REG,
	input logic [31:0] DMA1CNT_L_REG,
	input logic [31:0] DMA1CNT_H_REG,
	input logic [31:0] DMA2SAD_L_REG,
	input logic [31:0] DMA2SAD_H_REG,
	input logic [31:0] DMA2DAD_L_REG,
	input logic [31:0] DMA2DAD_H_REG,
	input logic [31:0] DMA2CNT_L_REG,
	input logic [31:0] DMA2CNT_H_REG,
	input logic [31:0] DMA3SAD_L_REG,
	input logic [31:0] DMA3SAD_H_REG,
	input logic [31:0] DMA3DAD_L_REG,
	input logic [31:0] DMA3DAD_H_REG,
	input logic [31:0] DMA3CNT_L_REG,
	input logic [31:0] DMA3CNT_H_REG,
   
   input  logic [15:0] vcount, hcount,
   input  logic cpu_preemptable,
   input  logic        sound_req1, sound_req2,

   input  logic        mem_wait,

   input  logic [31:0] rdata,
   output wire  [31:0] addr,
   output wire  [31:0] wdata,
   output wire  [1:0]  size,
   output wire         wen,

   output logic [3:0]  disable_dma,
   output logic        active,
   output logic        irq0, irq1, irq2, irq3,

   input  logic clk, rst_b);

   logic [15:0] controlL0, controlH0;
   logic [15:0] srcAddrL0, srcAddrH0;
   logic [15:0] destAddrL0, destAddrH0;

   logic [15:0] controlL1, controlH1;
   logic [15:0] srcAddrL1, srcAddrH1;
   logic [15:0] destAddrL1, destAddrH1;

   logic [15:0] controlL2, controlH2;
   logic [15:0] srcAddrL2, srcAddrH2;
   logic [15:0] destAddrL2, destAddrH2;

   logic [15:0] controlL3, controlH3;
   logic [15:0] srcAddrL3, srcAddrH3;
   logic [15:0] destAddrL3, destAddrH3;

   assign controlL0 = DMA0CNT_L_REG[15:0];
   assign controlH0 = DMA0CNT_H_REG[31:16];
   assign srcAddrL0 = DMA0SAD_L_REG[15:0];
   assign srcAddrH0 = DMA0SAD_H_REG[31:16];
   assign destAddrL0 = DMA0DAD_L_REG[15:0];
   assign destAddrH0 = DMA0DAD_H_REG[31:16];

   assign controlL1 = DMA1CNT_L_REG[15:0];
   assign controlH1 = DMA1CNT_H_REG[31:16];
   assign srcAddrL1 = DMA1SAD_L_REG[15:0];
   assign srcAddrH1 = DMA1SAD_H_REG[31:16];
   assign destAddrL1 = DMA1DAD_L_REG[15:0];
   assign destAddrH1 = DMA1DAD_H_REG[31:16];

   assign controlL2 = DMA2CNT_L_REG[15:0];
   assign controlH2 = DMA2CNT_H_REG[31:16];
   assign srcAddrL2 = DMA2SAD_L_REG[15:0];
   assign srcAddrH2 = DMA2SAD_H_REG[31:16];
   assign destAddrL2 = DMA2DAD_L_REG[15:0];
   assign destAddrH2 = DMA2DAD_H_REG[31:16];

   assign controlL3 = DMA3CNT_L_REG[15:0];
   assign controlH3 = DMA3CNT_H_REG[31:16];
   assign srcAddrL3 = DMA3SAD_L_REG[15:0];
   assign srcAddrH3 = DMA3SAD_H_REG[31:16];
   assign destAddrL3 = DMA3DAD_L_REG[15:0];
   assign destAddrH3 = DMA3DAD_H_REG[31:16];

   logic [3:0] preempts;
   (* mark_debug = "true" *) logic [3:0] actives;
   logic [3:0] mid_process;
   logic allowed_to_begin;

   assign active = |actives;
   assign preempts[0] = 1'b0;
   assign preempts[1] = actives[0];
   assign preempts[2] = actives[0] | actives[1];
   assign preempts[3] = actives[0] | actives[1] | actives[2];
   assign allowed_to_begin = ~mid_process[0] && ~mid_process[1]
                             && ~mid_process[2] && ~mid_process[3];


   dma_unit dma0(.controlL(controlL0), .controlH(controlH0),
                 .srcAddrL(srcAddrL0), .srcAddrH(srcAddrH0),
                 .destAddrL(destAddrL0), .destAddrH(destAddrH0),
                 .mem_wait, .preempted(preempts[0]),
                 .srcGamePak(1'b0), .destGamePak(1'b0),
                 .disable_dma(disable_dma[0]),
                 .active(actives[0]), .allowed_to_begin,
                 .irq(irq0), .others_cant_preempt(mid_process[0]),
                 .addr, .wdata, .rdata, .size, .wen,
                 .vcount, .hcount, .sound(1'b0), .sound_req(1'b0),
                 .cpu_preemptable,
                 .clk, .rst_b);

   dma_unit dma1(.controlL(controlL1), .controlH(controlH1),
                 .srcAddrL(srcAddrL1), .srcAddrH(srcAddrH1),
                 .destAddrL(destAddrL1), .destAddrH(destAddrH1),
                 .mem_wait, .preempted(preempts[1]),
                 .srcGamePak(1'b1), .destGamePak(1'b0),
                 .disable_dma(disable_dma[1]),
                 .active(actives[1]), .allowed_to_begin,
                 .irq(irq1), .others_cant_preempt(mid_process[1]),
                 .addr, .wdata, .rdata, .size, .wen,
                 .vcount, .hcount, .sound(1'b1), .sound_req(sound_req1),
                 .cpu_preemptable,
                 .clk, .rst_b);

   dma_unit dma2(.controlL(controlL2), .controlH(controlH2),
                 .srcAddrL(srcAddrL2), .srcAddrH(srcAddrH2),
                 .destAddrL(destAddrL2), .destAddrH(destAddrH2),
                 .mem_wait, .preempted(preempts[2]),
                 .srcGamePak(1'b1), .destGamePak(1'b0),
                 .disable_dma(disable_dma[2]),
                 .active(actives[2]), .allowed_to_begin,
                 .irq(irq2), .others_cant_preempt(mid_process[2]),
                 .addr, .wdata, .rdata, .size, .wen,
                 .vcount, .hcount, .sound(1'b1), .sound_req(sound_req2),
                 .cpu_preemptable,
                 .clk, .rst_b);

   dma_unit dma3(.controlL(controlL3), .controlH(controlH3),
                 .srcAddrL(srcAddrL3), .srcAddrH(srcAddrH3),
                 .destAddrL(destAddrL3), .destAddrH(destAddrH3),
                 .mem_wait, .preempted(preempts[3]),
                 .srcGamePak(1'b1), .destGamePak(1'b1),
                 .disable_dma(disable_dma[3]),
                 .active(actives[3]), .allowed_to_begin,
                 .irq(irq3), .others_cant_preempt(mid_process[3]),
                 .addr, .wdata, .rdata, .size, .wen,
                 .vcount, .hcount, .sound(1'b0), .sound_req(1'b0),
                 .cpu_preemptable,
                 .clk, .rst_b);

endmodule: dma_top

`default_nettype wire
